--background code when we learn sprites and shit