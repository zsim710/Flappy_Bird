--lives shit here