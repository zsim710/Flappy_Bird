--A graphical way of checking score using 7 segment display