--ground code for when the ground is needed